// This module contains a Verilog description of the top level module
// Assuming you don't modify the inputs and outputs of the various submodules,
// you should not have to modify anything in this file.

module task7(input CLOCK_50, input[3:0] KEY, output[9:0] LEDR,
            output[6:0] HEX5, output[6:0] HEX4, output[6:0] HEX3,
            output[6:0] HEX2, output[6:0] HEX1, output[6:0] HEX0
            /* any other signals you need */ );

endmodule

