module card7seg(input logic [3:0] SW, output logic [6:0] HEX0);
		
   // your code goes here
	
endmodule

