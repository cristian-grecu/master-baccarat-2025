module card7seg(input logic [3:0] card, output logic [6:0] seg7);

   // your code goes here

endmodule

